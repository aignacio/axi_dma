`ifndef _DMA_UTILS_PKG_
`define _DMA_UTILS_PKG_
  package dma_utils_pkg;
    //export *::*;
    `include "dma_axi_pkg.svh"
    `include "dma_pkg.svh"
  endpackage
`endif
