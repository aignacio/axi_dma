`ifndef _UTILS_PKG_
`define _UTILS_PKG_
  package utils_pkg;
    //export *::*;
    `include "axi_pkg.svh"
    `include "dma_pkg.svh"
  endpackage
`endif
