`ifndef _DMA_UTILS_PKG_
`define _DMA_UTILS_PKG_
  package dma_utils_pkg;
    `include "dma_pkg.svh"
  endpackage
`endif
